** Profile: "SCHEMATIC1-TEST"  [ D:\Otros\Electr�nica\PhonoPreamp\Simulations\phonopreamp-pspicefiles\schematic1\test.sim ] 

** Creating circuit file "TEST.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 20 20000
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
